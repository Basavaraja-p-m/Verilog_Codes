module encoder_8b10b (
    input  [7:0] data_in,   
    input  rd,
    input  k,
    output reg [9:0] data_out    
              );

always @(*) begin
   if (k) begin
       case (data_in)
    8'h1C: data_out = rd ? 10'b0011110100 : 10'b1100001011;
    8'h3C: data_out = rd ? 10'b0011111001 : 10'b1100000110;
    8'h5C: data_out = rd ? 10'b0011110101 : 10'b1100001010;
    8'h7C: data_out = rd ? 10'b0011110011 : 10'b1100001100;
    8'h9C: data_out = rd ? 10'b0011110010 : 10'b1100001101;

    8'hBC: data_out = rd ? 10'b0011111010 : 10'b1100000101;
    8'hDC: data_out = rd ? 10'b0011110110 : 10'b1100001001;
    8'hFC: data_out = rd ? 10'b0011111000 : 10'b1100000111;
    8'hF7: data_out = rd ? 10'b1110101000 : 10'b0001010111;
    8'hFB: data_out = rd ? 10'b1101101000 : 10'b0010010111;

    8'hFD: data_out = rd ? 10'b1011101000 : 10'b0100010111;
    8'hFE: data_out = rd ? 10'b0111101000 : 10'b1000010111;         
   endcase
 end
    else 
        begin
           case (data_in)

        8'h00: data_out = (rd) ? 10'b1001110100 : 10'b0110001011; 
        8'h01: data_out = (rd) ? 10'b0111010100 : 10'b1000101011; 
        8'h02: data_out = (rd) ? 10'b1011010100 : 10'b0100101011; 
        8'h03: data_out = (rd) ? 10'b1100011011 : 10'b1100010100; 
        8'h04: data_out = (rd) ? 10'b1101010100 : 10'b0010101011;
		
        8'h05: data_out = (rd) ? 10'b1010011011 : 10'b1010010100; 
        8'h06: data_out = (rd) ? 10'b0110011011 : 10'b0110010100; 
        8'h07: data_out = (rd) ? 10'b1110001011 : 10'b0001110100; 
        8'h08: data_out = (rd) ? 10'b1110010100 : 10'b0001101011; 
        8'h09: data_out = (rd) ? 10'b1001011011 : 10'b1001010100; 
		
        8'h0A: data_out = (rd) ? 10'b0101011011 : 10'b0101010100; 
        8'h0B: data_out = (rd) ? 10'b1101001011 : 10'b1101000100; 
        8'h0C: data_out = (rd) ? 10'b0011011011 : 10'b0011010100; 
        8'h0D: data_out = (rd) ? 10'b1011001011 : 10'b1011000100; 
        8'h0E: data_out = (rd) ? 10'b0111001011 : 10'b0111000100; 

        8'h0F: data_out = (rd) ? 10'b0101110100 : 10'b1010001011; 
        8'h10: data_out = rd ? 10'b0110110100 : 10'b1001001011;
    	8'h11: data_out = rd ? 10'b1000111011 : 10'b1000110100;
    	8'h12: data_out = rd ? 10'b0100111011 : 10'b0100110100;
   	 	8'h13: data_out = rd ? 10'b1100101011 : 10'b1100100100;

    	8'h14: data_out = rd ? 10'b0010111011 : 10'b0010110100;
   	 	8'h15: data_out = rd ? 10'b1010101011 : 10'b1010100100;
    	8'h16: data_out = rd ? 10'b0110101011 : 10'b0110100100;
    	8'h17: data_out = rd ? 10'b1110100100 : 10'b0001011011;
    	8'h18: data_out = rd ? 10'b1100110100 : 10'b0011001011;

    	8'h19: data_out = rd ? 10'b1001101011 : 10'b1001100100;
   		8'h1A: data_out = rd ? 10'b0101101011 : 10'b0101100100;
    	8'h1B: data_out = rd ? 10'b1101100100 : 10'b0010011011;
    	8'h1C: data_out = rd ? 10'b0011101011 : 10'b0011100100;
    	8'h1D: data_out = rd ? 10'b1011100100 : 10'b0100011011;
		
    8'h1E: data_out = rd ? 10'b0111100100 : 10'b1000011011;
    8'h1F: data_out = rd ? 10'b1010110100 : 10'b0101001011;
    8'h20: data_out = rd ? 10'b1001111001 : 10'b0110001001;
    8'h21: data_out = rd ? 10'b0111011001 : 10'b1000101001;
    8'h22: data_out = rd ? 10'b1011011001 : 10'b0100101001;

    8'h23: data_out = rd ? 10'b1100011001 : 10'b1100011001;
    8'h24: data_out = rd ? 10'b1101011001 : 10'b0010101001;
    8'h25: data_out = rd ? 10'b1010011001 : 10'b1010011001;
    8'h26: data_out = rd ? 10'b0110011001 : 10'b0110011001;
    8'h27: data_out = rd ? 10'b1110001001 : 10'b0001111001;
	
    8'h28: data_out = rd ? 10'b1110011001 : 10'b0001101001;
    8'h29: data_out = rd ? 10'b1001011001 : 10'b1001011001;
    8'h2A: data_out = rd ? 10'b0101011001 : 10'b0101011001;
    8'h2B: data_out = rd ? 10'b1101001001 : 10'b1101001001;
    8'h2C: data_out = rd ? 10'b0011011001 : 10'b0011011001;
    8'h2D: data_out = rd ? 10'b1011001001 : 10'b1011001001;

	8'h2E: data_out = rd ? 10'b0111001001 : 10'b0111001001;
    8'h2F: data_out = rd ? 10'b0101111001 : 10'b1010001001;
    8'h30: data_out = rd ? 10'b0110111001 : 10'b1001001001;
    8'h31: data_out = rd ? 10'b1000111001 : 10'b1000111001;
    8'h32: data_out = rd ? 10'b0100111001 : 10'b0100111001;

    8'h33: data_out = rd ? 10'b1100101001 : 10'b1100101001;
    8'h34: data_out = rd ? 10'b0010111001 : 10'b0010111001;
    8'h35: data_out = rd ? 10'b1010101001 : 10'b1010101001;
    8'h36: data_out = rd ? 10'b0110101001 : 10'b0110101001;
    8'h37: data_out = rd ? 10'b1110101001 : 10'b0001011001;

    8'h38: data_out = rd ? 10'b1100111001 : 10'b0011001001;
    8'h39: data_out = rd ? 10'b1001101001 : 10'b1001101001;
    8'h3A: data_out = rd ? 10'b0101101001 : 10'b0101101001;
    8'h3B: data_out = rd ? 10'b1101101001 : 10'b0010011001;
    8'h3C: data_out = rd ? 10'b0011101001 : 10'b0011101001;

    8'h3D: data_out = rd ? 10'b1011101001 : 10'b0100011001;
    8'h3E: data_out = rd ? 10'b0111101001 : 10'b1000011001;
    8'h3F: data_out = rd ? 10'b1010111001 : 10'b0101001001;
    8'h40: data_out = rd ? 10'b1001110101 : 10'b0110000101;
    8'h41: data_out = rd ? 10'b0111010101 : 10'b1000100101;

    8'h42: data_out = rd ? 10'b1011010101 : 10'b0100100101;
    8'h43: data_out = rd ? 10'b1100010101 : 10'b1100010101;
    8'h44: data_out = rd ? 10'b1101010101 : 10'b0010100101;
    8'h45: data_out = rd ? 10'b1010010101 : 10'b1010010101;
    8'h46: data_out = rd ? 10'b0110010101 : 10'b0110010101;

    8'h47: data_out = rd ? 10'b1110000101 : 10'b0001110101;
    8'h48: data_out = rd ? 10'b1110010101 : 10'b0001100101;
    8'h49: data_out = rd ? 10'b1001010101 : 10'b1001010101;
    8'h4A: data_out = rd ? 10'b0101010101 : 10'b0101010101;
    8'h4B: data_out = rd ? 10'b1101000101 : 10'b1101000101;

    8'h4C: data_out = rd ? 10'b0011010101 : 10'b0011010101;
    8'h4D: data_out = rd ? 10'b1011000101 : 10'b1011000101;
    8'h4E: data_out = rd ? 10'b0111000101 : 10'b0111000101;
    8'h4F: data_out = rd ? 10'b0101110101 : 10'b1010000101;
    8'h50: data_out = rd ? 10'b0110110101 : 10'b1001000101;

    8'h51: data_out = rd ? 10'b1000110101 : 10'b1000110101;
    8'h52: data_out = rd ? 10'b0100110101 : 10'b0100110101;
    8'h53: data_out = rd ? 10'b1100100101 : 10'b1100100101;
    8'h54: data_out = rd ? 10'b0010110101 : 10'b0010110101;
    8'h55: data_out = rd ? 10'b1010100101 : 10'b1010100101;

    8'h56: data_out = rd ? 10'b0110100101 : 10'b0110100101;
    8'h57: data_out = rd ? 10'b1110100101 : 10'b0001010101;
    8'h58: data_out = rd ? 10'b1100110101 : 10'b0011000101;
	
    8'h59: data_out = rd ? 10'b1001100101 : 10'b1001100101;
    8'h5A: data_out = rd ? 10'b0101100101 : 10'b0101100101;
    8'h5B: data_out = rd ? 10'b1101100101 : 10'b0010010101;
    8'h5C: data_out = rd ? 10'b0011100101 : 10'b0011100101;
    8'h5D: data_out = rd ? 10'b1011100101 : 10'b0100010101;

    8'h5E: data_out = rd ? 10'b0111100101 : 10'b1000010101;
    8'h5F: data_out = rd ? 10'b1010110101 : 10'b0101000101; 
    8'h60: data_out = rd ? 10'b1001110011 : 10'b0110001100;
    8'h61: data_out = rd ? 10'b0111010011 : 10'b1000101100;
    8'h62: data_out = rd ? 10'b1011010011 : 10'b0100101100;

    8'h63: data_out = rd ? 10'b1100011100 : 10'b1100010011;
    8'h64: data_out = rd ? 10'b1101010011 : 10'b0010101100;
    8'h65: data_out = rd ? 10'b1010011100 : 10'b1010010011;
    8'h66: data_out = rd ? 10'b0110011100 : 10'b0110010011;
    8'h67: data_out = rd ? 10'b1110001100 : 10'b0001110011;
	
    8'h68: data_out = rd ? 10'b1110010011 : 10'b0001101100;
    8'h69: data_out = rd ? 10'b1001011100 : 10'b1001010011;
    8'h6A: data_out = rd ? 10'b0101011100 : 10'b0101010011;
    8'h6B: data_out = rd ? 10'b1101001100 : 10'b110100011;
    8'h6C: data_out = rd ? 10'b0011011100 : 10'b0011010011;

    8'h6D: data_out = rd ? 10'b1011001100 : 10'b101100011;
    8'h6E: data_out = rd ? 10'b0111001100 : 10'b011100011;
    8'h6F: data_out = rd ? 10'b0101110011 : 10'b1010001100;
    8'h70: data_out = rd ? 10'b0110110011 : 10'b1001001100;
    8'h71: data_out = rd ? 10'b1000111100 : 10'b1000110011;

    8'h72: data_out = rd ? 10'b0100111100 : 10'b0100110011;
    8'h73: data_out = rd ? 10'b1100101100 : 10'b1100100011;
    8'h74: data_out = rd ? 10'b0010111100 : 10'b0010110011;
    8'h75: data_out = rd ? 10'b1010101100 : 10'b1010100011;
    8'h76: data_out = rd ? 10'b0110101100 : 10'b0110100011;

    8'h77: data_out = rd ? 10'b1110100011 : 10'b0001011100;
    8'h78: data_out = rd ? 10'b1100110011 : 10'b0011001100;
    8'h79: data_out = rd ? 10'b1001101100 : 10'b1001100011;
	
    8'h7A: data_out = rd ? 10'b0101101100 : 10'b0101100011;
    8'h7B: data_out = rd ? 10'b1101100011 : 10'b0010011100;
    8'h7C: data_out = rd ? 10'b0011101100 : 10'b0011100011;
    8'h7D: data_out = rd ? 10'b1011100011 : 10'b0100011100;
    8'h7E: data_out = rd ? 10'b0111100011 : 10'b1000011100;

    8'h7F: data_out = rd ? 10'b1010110011 : 10'b0101001100;
    8'h80: data_out = rd ? 10'b1001110010 : 10'b0110001101;
    8'h81: data_out = rd ? 10'b0111010010 : 10'b1000101101;
    8'h82: data_out = rd ? 10'b1011010010 : 10'b0100101101;
    8'h83: data_out = rd ? 10'b1100011101 : 10'b1100010010;

    8'h84: data_out = rd ? 10'b1101010010 : 10'b0010101101;
	8'h85: data_out = rd ? 10'b1010011101 : 10'b1010010010;
    8'h86: data_out = rd ? 10'b0110011101 : 10'b0110010010;
    8'h87: data_out = rd ? 10'b1110001101 : 10'b0001110010;
    8'h88: data_out = rd ? 10'b1110010010 : 10'b0001101101;

    8'h89: data_out = rd ? 10'b1001011101 : 10'b1001010010;
    8'h8A: data_out = rd ? 10'b0101011101 : 10'b0101010010;
    8'h8B: data_out = rd ? 10'b1101001101 : 10'b0010100010;
    8'h8C: data_out = rd ? 10'b0011011101 : 10'b0011010010;
    8'h8D: data_out = rd ? 10'b1011001101 : 10'b1011000010;

    8'h8E: data_out = rd ? 10'b0111001101 : 10'b0111000010;
    8'h8F: data_out = rd ? 10'b0101110010 : 10'b1010001101;
    8'h90: data_out = rd ? 10'b0110110010 : 10'b1001001101;
    8'h91: data_out = rd ? 10'b1000111101 : 10'b1000110010;
    8'h92: data_out = rd ? 10'b0100111101 : 10'b0100110010;

    8'h93: data_out = rd ? 10'b1100101101 : 10'b1100100010;
    8'h94: data_out = rd ? 10'b0010111101 : 10'b0010110010;
    8'h95: data_out = rd ? 10'b1010101101 : 10'b1010100010;
    8'h96: data_out = rd ? 10'b0110101101 : 10'b0110100010;
    8'h97: data_out = rd ? 10'b1110100010 : 10'b0001011101;

	8'h98: data_out = rd ? 10'b1100110010 : 10'b0011001101;
    8'h99: data_out = rd ? 10'b1001101101 : 10'b1001100010;
    8'h9A: data_out = rd ? 10'b0101101101 : 10'b0101100010;
	
    8'h9B: data_out = rd ? 10'b1101100010 : 10'b0010011101;
    8'h9C: data_out = rd ? 10'b0011101101 : 10'b0011100010;
    8'h9D: data_out = rd ? 10'b1011100010 : 10'b0100011101;
    8'h9E: data_out = rd ? 10'b0111100010 : 10'b1000011101;
    8'h9F: data_out = rd ? 10'b1010110010 : 10'b0101001101;
	
    8'hA0: data_out = rd ? 10'b1001111010 : 10'b0110001010;
    8'hA1: data_out = rd ? 10'b0111011010 : 10'b1000101010;
    8'hA2: data_out = rd ? 10'b1011011010 : 10'b0100101010;
    8'hA3: data_out = rd ? 10'b1100011010 : 10'b1100011010;
    8'hA4: data_out = rd ? 10'b1101011010 : 10'b0010101010;

    8'hA5: data_out = rd ? 10'b1010011010 : 10'b1010011010;
    8'hA6: data_out = rd ? 10'b0110011010 : 10'b0110011010;
    8'hA7: data_out = rd ? 10'b1110001010 : 10'b0001111010;
    8'hA8: data_out = rd ? 10'b1110011010 : 10'b0001101010;
    8'hA9: data_out = rd ? 10'b1001011010 : 10'b1001011010;

    8'hAA: data_out = rd ? 10'b0101011010 : 10'b0101011010;
    8'hAB: data_out = rd ? 10'b1101001010 : 10'b1101001010;
    8'hAC: data_out = rd ? 10'b0011011010 : 10'b0011011010;
    8'hAD: data_out = rd ? 10'b1011001010 : 10'b1011001010;
    8'hAE: data_out = rd ? 10'b0111001010 : 10'b0111001010;

    8'hAF: data_out = rd ? 10'b0101111010 : 10'b1010001010;
    8'hB0: data_out = rd ? 10'b0110111010 : 10'b1001001010;
    8'hB1: data_out = rd ? 10'b1000111010 : 10'b1000111010;
    8'hB2: data_out = rd ? 10'b0100111010 : 10'b0100111010;
    8'hB3: data_out = rd ? 10'b1100101010 : 10'b1100101010;

    8'hB4: data_out = rd ? 10'b0010111010 : 10'b0010111010;
    8'hB5: data_out = rd ? 10'b1010101010 : 10'b1010101010;
    8'hB6: data_out = rd ? 10'b0110101010 : 10'b0110101010;
    8'hB7: data_out = rd ? 10'b1110101010 : 10'b0001011010;
    8'hB8: data_out = rd ? 10'b1100111010 : 10'b0011001010;

    8'hB9: data_out = rd ? 10'b1001101010 : 10'b1001101010;
    8'hBA: data_out = rd ? 10'b0101101010 : 10'b0101101010;
    8'hBB: data_out = rd ? 10'b1101101010 : 10'b0010011010;

    8'hBC: data_out = rd ? 10'b0011101010 : 10'b0011101010;
    8'hBD: data_out = rd ? 10'b1011101010 : 10'b0100011010;
    8'hBE: data_out = rd ? 10'b0111101010 : 10'b1000011010;
    8'hBF: data_out = rd ? 10'b1010111010 : 10'b0101001010; 
    8'hC0: data_out = rd ? 10'b1001110110 : 10'b0110000110;

    8'hC1: data_out = rd ? 10'b0111010110 : 10'b1000100110;
    8'hC2: data_out = rd ? 10'b1011010110 : 10'b0100100110;
    8'hC3: data_out = rd ? 10'b1100010110 : 10'b1100010110;
    8'hC4: data_out = rd ? 10'b1101010110 : 10'b0010100110;
    8'hC5: data_out = rd ? 10'b1010010110 : 10'b1010010110;

    8'hC6: data_out = rd ? 10'b0110010110 : 10'b0110010110;
    8'hC7: data_out = rd ? 10'b1110000110 : 10'b0001110110;
    8'hC8: data_out = rd ? 10'b1110010110 : 10'b0001100110;
    8'hC9: data_out = rd ? 10'b1001010110 : 10'b1001010110;
    8'hCA: data_out = rd ? 10'b0101010110 : 10'b0101010110;

    8'hCB: data_out = rd ? 10'b1101000110 : 10'b1101000110;
    8'hCC: data_out = rd ? 10'b0011010110 : 10'b0011010110;
    8'hCD: data_out = rd ? 10'b1011000110 : 10'b1011000110;
    8'hCE: data_out = rd ? 10'b0111000110 : 10'b0111000110;
    8'hCF: data_out = rd ? 10'b0101110110 : 10'b1010000110;

    8'hD0: data_out = rd ? 10'b0110110110 : 10'b1001000110;
    8'hD1: data_out = rd ? 10'b1000110110 : 10'b1000110110;
    8'hD2: data_out = rd ? 10'b0100110110 : 10'b0100110110;
    8'hD3: data_out = rd ? 10'b1100100110 : 10'b1100100110;
    8'hD4: data_out = rd ? 10'b0010110110 : 10'b0010110110;

    8'hD5: data_out = rd ? 10'b1010100110 : 10'b1010100110;
    8'hD6: data_out = rd ? 10'b0110100110 : 10'b0110100110;
    8'hD7: data_out = rd ? 10'b1110100110 : 10'b0001010110;
    8'hD8: data_out = rd ? 10'b1100110110 : 10'b0011000110;
    8'hD9: data_out = rd ? 10'b1001100110 : 10'b1001100110;

    8'hDA: data_out = rd ? 10'b0101100110 : 10'b0101100110;
    8'hDB: data_out = rd ? 10'b1101100110 : 10'b0010010110;
    8'hDC: data_out = rd ? 10'b0011100110 : 10'b0011100110;

    8'hDD: data_out = rd ? 10'b1011100110 : 10'b0100010110;
    8'hDE: data_out = rd ? 10'b0111100110 : 10'b1000010110;
    8'hDF: data_out = rd ? 10'b1010110110 : 10'b0101000110;
    8'hE0: data_out = rd ? 10'b1001110001 : 10'b0110001110;
    8'hE1: data_out = rd ? 10'b0111010001 : 10'b1000101110;
	
    8'hE2: data_out = rd ? 10'b1011010001 : 10'b0100101110;
    8'hE3: data_out = rd ? 10'b1100011110 : 10'b1100010001;
    8'hE4: data_out = rd ? 10'b1101010001 : 10'b0010101110;
    8'hE5: data_out = rd ? 10'b1010011110 : 10'b1010010001;
    8'hE6: data_out = rd ? 10'b0110011110 : 10'b0110010001;
	
    8'hE7: data_out = rd ? 10'b1110001110 : 10'b0001110001;
    8'hE8: data_out = rd ? 10'b1110010001 : 10'b0001101110;
    8'hE9: data_out = rd ? 10'b1001011110 : 10'b1001010001;
    8'hEA: data_out = rd ? 10'b0101011110 : 10'b0101010001;
    8'hEB: data_out = rd ? 10'b1101001110 : 10'b1101001000;
	
    8'hEC: data_out = rd ? 10'b0011011110 : 10'b0011010001;
    8'hED: data_out = rd ? 10'b1011001110 : 10'b1011001000;
    8'hEE: data_out = rd ? 10'b0111001110 : 10'b0111001000;
    8'hEF: data_out = rd ? 10'b0101110001 : 10'b1010001110;
    8'hF0: data_out = rd ? 10'b0110110001 : 10'b1001001110;
	
    8'hF1: data_out = rd ? 10'b1000110111 : 10'b1000110001;
    8'hF2: data_out = rd ? 10'b0100110111 : 10'b0100110001;
    8'hF3: data_out = rd ? 10'b1100101110 : 10'b1100100001;
    8'hF4: data_out = rd ? 10'b0010110111 : 10'b0010110001;
    8'hF5: data_out = rd ? 10'b1010101110 : 10'b1010100001;
	
    8'hF6: data_out = rd ? 10'b0110101110 : 10'b0110100001;
    8'hF7: data_out = rd ? 10'b1110100001 : 10'b0001011110;
    8'hF8: data_out = rd ? 10'b1100110001 : 10'b0011001110;
    8'hF9: data_out = rd ? 10'b1001101110 : 10'b1001100001;
    8'hFA: data_out = rd ? 10'b0101101110 : 10'b0101100001;
	
    8'hFB: data_out = rd ? 10'b1101100001 : 10'b0010011110;
    8'hFC: data_out = rd ? 10'b0011101110 : 10'b0011100001;
    8'hFD: data_out = rd ? 10'b1011100001 : 10'b0100011110;
	
    8'hFE: data_out = rd ? 10'b0111100001 : 10'b1000011110;
    8'hFF: data_out = rd ? 10'b1010110001 : 10'b0101001110;

    default: data_out = 10'b0000000000;

  endcase
end

//rd_next = ~rd;
end

endmodule

