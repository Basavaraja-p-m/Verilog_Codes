module snippet();

reg [7:0]mem[31:0][31:0];

endmodule
