module DT();
    reg a;
    wire b;
    tri1 c;
    tri0 d;
    wor e;
    wand f;
    supply1 g;
    supply0 h;
    tri i;
    integer j;
    real k;
    initial
    $display("a=%b b=%b c=%b d=%b e=%b f=%b g=%b h=%b i=%b j=%b k=%b",a,b,c,d,e,f,g,e,f,g,h);
 endmodule


