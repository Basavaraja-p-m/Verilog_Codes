module data_types();
    reg a;
    wire b;
    wor c;
    wand d;
    supply1 e;
    supply0 f;
    tri g;
    tri1 h;
    tri0 i;
    tri1 j;
    integer k;
    real l;
  initial 
   $display("a=%b b=%b c=%b d=%b e=%b f=%b g=%b h=%b i=%b j=%b k=%b l=%b",a,b,c,d,e,f,g,h,i,j,k,l);
endmodule
